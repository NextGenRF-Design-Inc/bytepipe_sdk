`timescale 1ps/1ps

module system_top (
  
  output  wire          adrv9001_csn,
  output  wire          adrv9001_sclk,
  inout   wire          adrv9001_mosi,
  input   wire          adrv9001_miso,

  input  wire           adrv9001_dev_clk_in,
  output wire           adrv9001_rstn,
  output wire           adrv9001_tx1_en,
  output wire           adrv9001_tx2_en,
  output wire           adrv9001_rx1_en,
  output wire           adrv9001_rx2_en,
  input  wire           adrv9001_irq,
  inout  wire [11:0]    adrv9001_dgpio,  
  
  input  wire           adrv9001_rx1_dclk_n,
  input  wire           adrv9001_rx1_dclk_p,
  input  wire           adrv9001_rx1_idata_n,
  input  wire           adrv9001_rx1_idata_p,
  input  wire           adrv9001_rx1_qdata_n,
  input  wire           adrv9001_rx1_qdata_p,
  input  wire           adrv9001_rx1_strobe_n,
  input  wire           adrv9001_rx1_strobe_p,

  input  wire           adrv9001_rx2_dclk_n,
  input  wire           adrv9001_rx2_dclk_p,
  input  wire           adrv9001_rx2_idata_n,
  input  wire           adrv9001_rx2_idata_p,
  input  wire           adrv9001_rx2_qdata_n,
  input  wire           adrv9001_rx2_qdata_p,
  input  wire           adrv9001_rx2_strobe_n,
  input  wire           adrv9001_rx2_strobe_p,

  output wire           adrv9001_tx1_dclk_n,
  output wire           adrv9001_tx1_dclk_p,
  input  wire           adrv9001_tx1_ref_clk_n,
  input  wire           adrv9001_tx1_ref_clk_p,
  output wire           adrv9001_tx1_idata_n,
  output wire           adrv9001_tx1_idata_p,
  output wire           adrv9001_tx1_qdata_n,
  output wire           adrv9001_tx1_qdata_p,
  output wire           adrv9001_tx1_strobe_n,
  output wire           adrv9001_tx1_strobe_p,
  
  output wire           adrv9001_tx2_dclk_n,
  output wire           adrv9001_tx2_dclk_p,
  input  wire           adrv9001_tx2_ref_clk_n,
  input  wire           adrv9001_tx2_ref_clk_p,
  output wire           adrv9001_tx2_idata_n,
  output wire           adrv9001_tx2_idata_p,
  output wire           adrv9001_tx2_qdata_n,
  output wire           adrv9001_tx2_qdata_p,
  output wire           adrv9001_tx2_strobe_n,
  output wire           adrv9001_tx2_strobe_p,
  input  wire  [ 3:0]   gpio_sw,
  input  wire  [ 2:0]   gpio_pb,
  output wire  [ 5:0]   gpio_led);
  
  system i_system (
    .dio_dev_clk                        (adrv9001_dev_clk_in),
    .dio_dgpio                          (adrv9001_dgpio),
    .dio_gp_int                         (adrv9001_irq),
    .dio_mode                           (),
    .dio_resetb                         (adrv9001_rstn),
    
    .dio_rx0_cssi_clk_lssi_clk_p        (adrv9001_rx1_dclk_p),
    .dio_rx0_cssi_data0_lssi_data0_n    (adrv9001_rx1_idata_n),
    .dio_rx0_cssi_data1_lssi_data0_p    (adrv9001_rx1_idata_p),
    .dio_rx0_cssi_data2_lssi_data1_n    (adrv9001_rx1_qdata_n),
    .dio_rx0_cssi_data3_lssi_data1_p    (adrv9001_rx1_qdata_p),
    .dio_rx0_cssi_gpio_enb              (),
    .dio_rx0_cssi_gpio_in               (8'd0),
    .dio_rx0_cssi_gpio_out              (),
    .dio_rx0_cssi_nc_lssi_clk_n         (adrv9001_rx1_dclk_n),
    .dio_rx0_cssi_nc_lssi_strobe_n      (adrv9001_rx1_strobe_n),
    .dio_rx0_cssi_strobe_lssi_strobe_p  (adrv9001_rx1_strobe_p),
    .dio_rx0_enable                     (adrv9001_rx1_en),
    
    .dio_rx1_cssi_clk_lssi_clk_p        (adrv9001_rx2_dclk_p),
    .dio_rx1_cssi_data0_lssi_data0_n    (adrv9001_rx2_idata_n),
    .dio_rx1_cssi_data1_lssi_data0_p    (adrv9001_rx2_idata_p),
    .dio_rx1_cssi_data2_lssi_data1_n    (adrv9001_rx2_qdata_n),
    .dio_rx1_cssi_data3_lssi_data1_p    (adrv9001_rx2_qdata_p),
    .dio_rx1_cssi_gpio_enb              (),
    .dio_rx1_cssi_gpio_in               (8'd0),
    .dio_rx1_cssi_gpio_out              (),
    .dio_rx1_cssi_nc_lssi_clk_n         (adrv9001_rx2_dclk_n),
    .dio_rx1_cssi_nc_lssi_strobe_n      (adrv9001_rx2_strobe_n),
    .dio_rx1_cssi_strobe_lssi_strobe_p  (adrv9001_rx2_strobe_p),
    .dio_rx1_enable                     (adrv9001_rx2_en),
    
    .dio_tx0_cssi_clk_lssi_clk_p        (adrv9001_tx1_dclk_p),
    .dio_tx0_cssi_data0_lssi_data0_n    (adrv9001_tx1_idata_n),
    .dio_tx0_cssi_data1_lssi_data0_p    (adrv9001_tx1_idata_p),
    .dio_tx0_cssi_data2_lssi_data1_n    (adrv9001_tx1_qdata_n),
    .dio_tx0_cssi_data3_lssi_data1_p    (adrv9001_tx1_qdata_p),
    .dio_tx0_cssi_gpio_enb              (),
    .dio_tx0_cssi_gpio_in               (10'd0),
    .dio_tx0_cssi_gpio_out              (),
    .dio_tx0_cssi_nc_lssi_clk_n         (adrv9001_tx1_dclk_n),
    .dio_tx0_cssi_nc_lssi_refclk_n      (adrv9001_tx1_ref_clk_n),
    .dio_tx0_cssi_nc_lssi_strobe_n      (adrv9001_tx1_strobe_n),
    .dio_tx0_cssi_refclk_lssi_refclk_p  (adrv9001_tx1_ref_clk_p),
    .dio_tx0_cssi_strobe_lssi_strobe_p  (adrv9001_tx1_strobe_p),
    .dio_tx0_enable                     (adrv9001_tx1_en),
    
    .dio_tx1_cssi_clk_lssi_clk_p        (adrv9001_tx2_dclk_p),
    .dio_tx1_cssi_data0_lssi_data0_n    (adrv9001_tx2_idata_n),
    .dio_tx1_cssi_data1_lssi_data0_p    (adrv9001_tx2_idata_p),
    .dio_tx1_cssi_data2_lssi_data1_n    (adrv9001_tx2_qdata_n),
    .dio_tx1_cssi_data3_lssi_data1_p    (adrv9001_tx2_qdata_p),
    .dio_tx1_cssi_gpio_enb              (),
    .dio_tx1_cssi_gpio_in               (10'd0),
    .dio_tx1_cssi_gpio_out              (),
    .dio_tx1_cssi_nc_lssi_clk_n         (adrv9001_tx2_dclk_n),
    .dio_tx1_cssi_nc_lssi_refclk_n      (adrv9001_tx2_ref_clk_n),
    .dio_tx1_cssi_nc_lssi_strobe_n      (adrv9001_tx2_strobe_n),
    .dio_tx1_cssi_refclk_lssi_refclk_p  (adrv9001_tx2_ref_clk_p),
    .dio_tx1_cssi_strobe_lssi_strobe_p  (adrv9001_tx2_strobe_p),
    .dio_tx1_enable                     (adrv9001_tx2_en),
    .spi_sclk                           (adrv9001_sclk),
    .spi_ssn                            (adrv9001_csn),
    .spi_miso                           (adrv9001_miso),
    .spi_mosi                           (adrv9001_mosi),
    .gpio_in                            ({gpio_pb, gpio_sw}),
    .gpio_out                           (gpio_led));
    

    

endmodule

// **********************************************************************************
// **********************************************************************************
